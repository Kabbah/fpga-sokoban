library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PushBoxMap is
	generic (
		MAP_WIDTH_BITS  : natural := 4;
		MAP_HEIGHT_BITS : natural := 4
	);
	port (
		display_x         : in unsigned(3 downto 0);
		display_y         : in unsigned(3 downto 0);
		display_pos_value : out unsigned(2 downto 0)
	);
end entity;

architecture archPushBoxMap of PushBoxMap is

-- Matriz do mapa
-- Bit 2: indica se é um objetivo ou não
-- Bits 1 downto 0: indica o que está no local:
--   00: Parede
--   01: Chão
--   10: Jogador
--   11: Caixa
type map_matrix_t is array(2**MAP_WIDTH_BITS-1 downto 0, 2**MAP_HEIGHT_BITS-1 downto 0) of unsigned(2 downto 0);
constant map_matrix : map_matrix_t := (("000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011"),
                                       ("100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111"),
                                       ("111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100"),
                                       ("011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000"),
                                       ("000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011"),
                                       ("100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111"),
                                       ("111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100"),
                                       ("011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000"),
                                       ("000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011"),
                                       ("100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111"),
                                       ("111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100"),
                                       ("011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000"),
                                       ("000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011", "000", "001", "010", "011"),
                                       ("100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111", "100", "101", "110", "111"),
                                       ("111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100", "111", "110", "101", "100"),
                                       ("011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000", "011", "010", "001", "000"));

begin
	display_pos_value <= map_matrix(to_integer(display_y), to_integer(display_x));
end architecture;
